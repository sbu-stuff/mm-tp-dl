*Auto-gererated 10-cell delay line circuit

V1 1 0 PULSE(0 1 0 7.5n 7.5n 100n 1 1)
R1 1 0 220
C2 1 0 6.8p Cpar = 0
L2 1 2 290n
R3 2 3 0.17
C3 3 0 6.8p Cpar = 0
L3 3 4 290n
R4 4 5 0.17
C4 5 0 6.8p Cpar = 0
L4 5 6 290n
R5 6 7 0.17
C5 7 0 6.8p Cpar = 0
L5 7 8 290n
R6 8 9 0.17
C6 9 0 6.8p Cpar = 0
L6 9 10 290n
R7 10 11 0.17
C7 11 0 6.8p Cpar = 0
L7 11 12 290n
R8 12 13 0.17
C8 13 0 6.8p Cpar = 0
L8 13 14 290n
R9 14 15 0.17
C9 15 0 6.8p Cpar = 0
L9 15 16 290n
R10 16 17 0.17
C10 17 0 6.8p Cpar = 0
L10 17 18 290n
R11 18 19 0.17
C11 19 0 6.8p Cpar = 0
L11 19 20 290n
R12 20 -1 0.17
C12 -1 0 6.8p Cpar = 0
R13 -1 0 220

.tran 216n